LIBRARY IEEE;
USE ieeee.std_logic_1164.all/

ENTITY schematic2 IS 
    PORT (
        a: IN STD_LOGIC;
        b: IN STD_LOGIC;
        c: IN STD_LOGIC;
        d, e: IN STD_LOGIC;
    );
END schematic2;

ARCHITECTURE behaviour OF schematic2 IS 
BEGIN 

END behaviour;